library verilog;
use verilog.vl_types.all;
entity ProcTest is
end ProcTest;
