module Stage1();
    input clk;
